magic
tech sky130A
magscale 1 2
timestamp 1635439965
<< obsli1 >>
rect 1104 2159 298816 177361
<< obsm1 >>
rect 290 1708 299722 177540
<< metal2 >>
rect 1306 179200 1362 180000
rect 3882 179200 3938 180000
rect 6550 179200 6606 180000
rect 9126 179200 9182 180000
rect 11794 179200 11850 180000
rect 14462 179200 14518 180000
rect 17038 179200 17094 180000
rect 19706 179200 19762 180000
rect 22282 179200 22338 180000
rect 24950 179200 25006 180000
rect 27618 179200 27674 180000
rect 30194 179200 30250 180000
rect 32862 179200 32918 180000
rect 35438 179200 35494 180000
rect 38106 179200 38162 180000
rect 40774 179200 40830 180000
rect 43350 179200 43406 180000
rect 46018 179200 46074 180000
rect 48594 179200 48650 180000
rect 51262 179200 51318 180000
rect 53930 179200 53986 180000
rect 56506 179200 56562 180000
rect 59174 179200 59230 180000
rect 61750 179200 61806 180000
rect 64418 179200 64474 180000
rect 67086 179200 67142 180000
rect 69662 179200 69718 180000
rect 72330 179200 72386 180000
rect 74906 179200 74962 180000
rect 77574 179200 77630 180000
rect 80242 179200 80298 180000
rect 82818 179200 82874 180000
rect 85486 179200 85542 180000
rect 88062 179200 88118 180000
rect 90730 179200 90786 180000
rect 93398 179200 93454 180000
rect 95974 179200 96030 180000
rect 98642 179200 98698 180000
rect 101310 179200 101366 180000
rect 103886 179200 103942 180000
rect 106554 179200 106610 180000
rect 109130 179200 109186 180000
rect 111798 179200 111854 180000
rect 114466 179200 114522 180000
rect 117042 179200 117098 180000
rect 119710 179200 119766 180000
rect 122286 179200 122342 180000
rect 124954 179200 125010 180000
rect 127622 179200 127678 180000
rect 130198 179200 130254 180000
rect 132866 179200 132922 180000
rect 135442 179200 135498 180000
rect 138110 179200 138166 180000
rect 140778 179200 140834 180000
rect 143354 179200 143410 180000
rect 146022 179200 146078 180000
rect 148598 179200 148654 180000
rect 151266 179200 151322 180000
rect 153934 179200 153990 180000
rect 156510 179200 156566 180000
rect 159178 179200 159234 180000
rect 161754 179200 161810 180000
rect 164422 179200 164478 180000
rect 167090 179200 167146 180000
rect 169666 179200 169722 180000
rect 172334 179200 172390 180000
rect 174910 179200 174966 180000
rect 177578 179200 177634 180000
rect 180246 179200 180302 180000
rect 182822 179200 182878 180000
rect 185490 179200 185546 180000
rect 188066 179200 188122 180000
rect 190734 179200 190790 180000
rect 193402 179200 193458 180000
rect 195978 179200 196034 180000
rect 198646 179200 198702 180000
rect 201314 179200 201370 180000
rect 203890 179200 203946 180000
rect 206558 179200 206614 180000
rect 209134 179200 209190 180000
rect 211802 179200 211858 180000
rect 214470 179200 214526 180000
rect 217046 179200 217102 180000
rect 219714 179200 219770 180000
rect 222290 179200 222346 180000
rect 224958 179200 225014 180000
rect 227626 179200 227682 180000
rect 230202 179200 230258 180000
rect 232870 179200 232926 180000
rect 235446 179200 235502 180000
rect 238114 179200 238170 180000
rect 240782 179200 240838 180000
rect 243358 179200 243414 180000
rect 246026 179200 246082 180000
rect 248602 179200 248658 180000
rect 251270 179200 251326 180000
rect 253938 179200 253994 180000
rect 256514 179200 256570 180000
rect 259182 179200 259238 180000
rect 261758 179200 261814 180000
rect 264426 179200 264482 180000
rect 267094 179200 267150 180000
rect 269670 179200 269726 180000
rect 272338 179200 272394 180000
rect 274914 179200 274970 180000
rect 277582 179200 277638 180000
rect 280250 179200 280306 180000
rect 282826 179200 282882 180000
rect 285494 179200 285550 180000
rect 288070 179200 288126 180000
rect 290738 179200 290794 180000
rect 293406 179200 293462 180000
rect 295982 179200 296038 180000
rect 298650 179200 298706 180000
rect 294 0 350 800
rect 846 0 902 800
rect 1490 0 1546 800
rect 2042 0 2098 800
rect 2686 0 2742 800
rect 3330 0 3386 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5722 0 5778 800
rect 6366 0 6422 800
rect 6918 0 6974 800
rect 7562 0 7618 800
rect 8114 0 8170 800
rect 8758 0 8814 800
rect 9402 0 9458 800
rect 9954 0 10010 800
rect 10598 0 10654 800
rect 11242 0 11298 800
rect 11794 0 11850 800
rect 12438 0 12494 800
rect 12990 0 13046 800
rect 13634 0 13690 800
rect 14278 0 14334 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16026 0 16082 800
rect 16670 0 16726 800
rect 17314 0 17370 800
rect 17866 0 17922 800
rect 18510 0 18566 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20350 0 20406 800
rect 20902 0 20958 800
rect 21546 0 21602 800
rect 22190 0 22246 800
rect 22742 0 22798 800
rect 23386 0 23442 800
rect 23938 0 23994 800
rect 24582 0 24638 800
rect 25226 0 25282 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27618 0 27674 800
rect 28262 0 28318 800
rect 28814 0 28870 800
rect 29458 0 29514 800
rect 30102 0 30158 800
rect 30654 0 30710 800
rect 31298 0 31354 800
rect 31850 0 31906 800
rect 32494 0 32550 800
rect 33138 0 33194 800
rect 33690 0 33746 800
rect 34334 0 34390 800
rect 34978 0 35034 800
rect 35530 0 35586 800
rect 36174 0 36230 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38566 0 38622 800
rect 39210 0 39266 800
rect 39762 0 39818 800
rect 40406 0 40462 800
rect 41050 0 41106 800
rect 41602 0 41658 800
rect 42246 0 42302 800
rect 42890 0 42946 800
rect 43442 0 43498 800
rect 44086 0 44142 800
rect 44638 0 44694 800
rect 45282 0 45338 800
rect 45926 0 45982 800
rect 46478 0 46534 800
rect 47122 0 47178 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49514 0 49570 800
rect 50158 0 50214 800
rect 50802 0 50858 800
rect 51354 0 51410 800
rect 51998 0 52054 800
rect 52550 0 52606 800
rect 53194 0 53250 800
rect 53838 0 53894 800
rect 54390 0 54446 800
rect 55034 0 55090 800
rect 55586 0 55642 800
rect 56230 0 56286 800
rect 56874 0 56930 800
rect 57426 0 57482 800
rect 58070 0 58126 800
rect 58714 0 58770 800
rect 59266 0 59322 800
rect 59910 0 59966 800
rect 60462 0 60518 800
rect 61106 0 61162 800
rect 61750 0 61806 800
rect 62302 0 62358 800
rect 62946 0 63002 800
rect 63498 0 63554 800
rect 64142 0 64198 800
rect 64786 0 64842 800
rect 65338 0 65394 800
rect 65982 0 66038 800
rect 66534 0 66590 800
rect 67178 0 67234 800
rect 67822 0 67878 800
rect 68374 0 68430 800
rect 69018 0 69074 800
rect 69662 0 69718 800
rect 70214 0 70270 800
rect 70858 0 70914 800
rect 71410 0 71466 800
rect 72054 0 72110 800
rect 72698 0 72754 800
rect 73250 0 73306 800
rect 73894 0 73950 800
rect 74446 0 74502 800
rect 75090 0 75146 800
rect 75734 0 75790 800
rect 76286 0 76342 800
rect 76930 0 76986 800
rect 77574 0 77630 800
rect 78126 0 78182 800
rect 78770 0 78826 800
rect 79322 0 79378 800
rect 79966 0 80022 800
rect 80610 0 80666 800
rect 81162 0 81218 800
rect 81806 0 81862 800
rect 82358 0 82414 800
rect 83002 0 83058 800
rect 83646 0 83702 800
rect 84198 0 84254 800
rect 84842 0 84898 800
rect 85486 0 85542 800
rect 86038 0 86094 800
rect 86682 0 86738 800
rect 87234 0 87290 800
rect 87878 0 87934 800
rect 88522 0 88578 800
rect 89074 0 89130 800
rect 89718 0 89774 800
rect 90270 0 90326 800
rect 90914 0 90970 800
rect 91558 0 91614 800
rect 92110 0 92166 800
rect 92754 0 92810 800
rect 93398 0 93454 800
rect 93950 0 94006 800
rect 94594 0 94650 800
rect 95146 0 95202 800
rect 95790 0 95846 800
rect 96434 0 96490 800
rect 96986 0 97042 800
rect 97630 0 97686 800
rect 98182 0 98238 800
rect 98826 0 98882 800
rect 99470 0 99526 800
rect 100022 0 100078 800
rect 100666 0 100722 800
rect 101310 0 101366 800
rect 101862 0 101918 800
rect 102506 0 102562 800
rect 103058 0 103114 800
rect 103702 0 103758 800
rect 104346 0 104402 800
rect 104898 0 104954 800
rect 105542 0 105598 800
rect 106094 0 106150 800
rect 106738 0 106794 800
rect 107382 0 107438 800
rect 107934 0 107990 800
rect 108578 0 108634 800
rect 109222 0 109278 800
rect 109774 0 109830 800
rect 110418 0 110474 800
rect 110970 0 111026 800
rect 111614 0 111670 800
rect 112258 0 112314 800
rect 112810 0 112866 800
rect 113454 0 113510 800
rect 114006 0 114062 800
rect 114650 0 114706 800
rect 115294 0 115350 800
rect 115846 0 115902 800
rect 116490 0 116546 800
rect 117134 0 117190 800
rect 117686 0 117742 800
rect 118330 0 118386 800
rect 118882 0 118938 800
rect 119526 0 119582 800
rect 120170 0 120226 800
rect 120722 0 120778 800
rect 121366 0 121422 800
rect 121918 0 121974 800
rect 122562 0 122618 800
rect 123206 0 123262 800
rect 123758 0 123814 800
rect 124402 0 124458 800
rect 124954 0 125010 800
rect 125598 0 125654 800
rect 126242 0 126298 800
rect 126794 0 126850 800
rect 127438 0 127494 800
rect 128082 0 128138 800
rect 128634 0 128690 800
rect 129278 0 129334 800
rect 129830 0 129886 800
rect 130474 0 130530 800
rect 131118 0 131174 800
rect 131670 0 131726 800
rect 132314 0 132370 800
rect 132866 0 132922 800
rect 133510 0 133566 800
rect 134154 0 134210 800
rect 134706 0 134762 800
rect 135350 0 135406 800
rect 135994 0 136050 800
rect 136546 0 136602 800
rect 137190 0 137246 800
rect 137742 0 137798 800
rect 138386 0 138442 800
rect 139030 0 139086 800
rect 139582 0 139638 800
rect 140226 0 140282 800
rect 140778 0 140834 800
rect 141422 0 141478 800
rect 142066 0 142122 800
rect 142618 0 142674 800
rect 143262 0 143318 800
rect 143906 0 143962 800
rect 144458 0 144514 800
rect 145102 0 145158 800
rect 145654 0 145710 800
rect 146298 0 146354 800
rect 146942 0 146998 800
rect 147494 0 147550 800
rect 148138 0 148194 800
rect 148690 0 148746 800
rect 149334 0 149390 800
rect 149978 0 150034 800
rect 150530 0 150586 800
rect 151174 0 151230 800
rect 151818 0 151874 800
rect 152370 0 152426 800
rect 153014 0 153070 800
rect 153566 0 153622 800
rect 154210 0 154266 800
rect 154854 0 154910 800
rect 155406 0 155462 800
rect 156050 0 156106 800
rect 156602 0 156658 800
rect 157246 0 157302 800
rect 157890 0 157946 800
rect 158442 0 158498 800
rect 159086 0 159142 800
rect 159730 0 159786 800
rect 160282 0 160338 800
rect 160926 0 160982 800
rect 161478 0 161534 800
rect 162122 0 162178 800
rect 162766 0 162822 800
rect 163318 0 163374 800
rect 163962 0 164018 800
rect 164514 0 164570 800
rect 165158 0 165214 800
rect 165802 0 165858 800
rect 166354 0 166410 800
rect 166998 0 167054 800
rect 167642 0 167698 800
rect 168194 0 168250 800
rect 168838 0 168894 800
rect 169390 0 169446 800
rect 170034 0 170090 800
rect 170678 0 170734 800
rect 171230 0 171286 800
rect 171874 0 171930 800
rect 172426 0 172482 800
rect 173070 0 173126 800
rect 173714 0 173770 800
rect 174266 0 174322 800
rect 174910 0 174966 800
rect 175554 0 175610 800
rect 176106 0 176162 800
rect 176750 0 176806 800
rect 177302 0 177358 800
rect 177946 0 178002 800
rect 178590 0 178646 800
rect 179142 0 179198 800
rect 179786 0 179842 800
rect 180338 0 180394 800
rect 180982 0 181038 800
rect 181626 0 181682 800
rect 182178 0 182234 800
rect 182822 0 182878 800
rect 183374 0 183430 800
rect 184018 0 184074 800
rect 184662 0 184718 800
rect 185214 0 185270 800
rect 185858 0 185914 800
rect 186502 0 186558 800
rect 187054 0 187110 800
rect 187698 0 187754 800
rect 188250 0 188306 800
rect 188894 0 188950 800
rect 189538 0 189594 800
rect 190090 0 190146 800
rect 190734 0 190790 800
rect 191286 0 191342 800
rect 191930 0 191986 800
rect 192574 0 192630 800
rect 193126 0 193182 800
rect 193770 0 193826 800
rect 194414 0 194470 800
rect 194966 0 195022 800
rect 195610 0 195666 800
rect 196162 0 196218 800
rect 196806 0 196862 800
rect 197450 0 197506 800
rect 198002 0 198058 800
rect 198646 0 198702 800
rect 199198 0 199254 800
rect 199842 0 199898 800
rect 200486 0 200542 800
rect 201038 0 201094 800
rect 201682 0 201738 800
rect 202326 0 202382 800
rect 202878 0 202934 800
rect 203522 0 203578 800
rect 204074 0 204130 800
rect 204718 0 204774 800
rect 205362 0 205418 800
rect 205914 0 205970 800
rect 206558 0 206614 800
rect 207110 0 207166 800
rect 207754 0 207810 800
rect 208398 0 208454 800
rect 208950 0 209006 800
rect 209594 0 209650 800
rect 210238 0 210294 800
rect 210790 0 210846 800
rect 211434 0 211490 800
rect 211986 0 212042 800
rect 212630 0 212686 800
rect 213274 0 213330 800
rect 213826 0 213882 800
rect 214470 0 214526 800
rect 215022 0 215078 800
rect 215666 0 215722 800
rect 216310 0 216366 800
rect 216862 0 216918 800
rect 217506 0 217562 800
rect 218150 0 218206 800
rect 218702 0 218758 800
rect 219346 0 219402 800
rect 219898 0 219954 800
rect 220542 0 220598 800
rect 221186 0 221242 800
rect 221738 0 221794 800
rect 222382 0 222438 800
rect 222934 0 222990 800
rect 223578 0 223634 800
rect 224222 0 224278 800
rect 224774 0 224830 800
rect 225418 0 225474 800
rect 226062 0 226118 800
rect 226614 0 226670 800
rect 227258 0 227314 800
rect 227810 0 227866 800
rect 228454 0 228510 800
rect 229098 0 229154 800
rect 229650 0 229706 800
rect 230294 0 230350 800
rect 230846 0 230902 800
rect 231490 0 231546 800
rect 232134 0 232190 800
rect 232686 0 232742 800
rect 233330 0 233386 800
rect 233974 0 234030 800
rect 234526 0 234582 800
rect 235170 0 235226 800
rect 235722 0 235778 800
rect 236366 0 236422 800
rect 237010 0 237066 800
rect 237562 0 237618 800
rect 238206 0 238262 800
rect 238758 0 238814 800
rect 239402 0 239458 800
rect 240046 0 240102 800
rect 240598 0 240654 800
rect 241242 0 241298 800
rect 241794 0 241850 800
rect 242438 0 242494 800
rect 243082 0 243138 800
rect 243634 0 243690 800
rect 244278 0 244334 800
rect 244922 0 244978 800
rect 245474 0 245530 800
rect 246118 0 246174 800
rect 246670 0 246726 800
rect 247314 0 247370 800
rect 247958 0 248014 800
rect 248510 0 248566 800
rect 249154 0 249210 800
rect 249706 0 249762 800
rect 250350 0 250406 800
rect 250994 0 251050 800
rect 251546 0 251602 800
rect 252190 0 252246 800
rect 252834 0 252890 800
rect 253386 0 253442 800
rect 254030 0 254086 800
rect 254582 0 254638 800
rect 255226 0 255282 800
rect 255870 0 255926 800
rect 256422 0 256478 800
rect 257066 0 257122 800
rect 257618 0 257674 800
rect 258262 0 258318 800
rect 258906 0 258962 800
rect 259458 0 259514 800
rect 260102 0 260158 800
rect 260746 0 260802 800
rect 261298 0 261354 800
rect 261942 0 261998 800
rect 262494 0 262550 800
rect 263138 0 263194 800
rect 263782 0 263838 800
rect 264334 0 264390 800
rect 264978 0 265034 800
rect 265530 0 265586 800
rect 266174 0 266230 800
rect 266818 0 266874 800
rect 267370 0 267426 800
rect 268014 0 268070 800
rect 268658 0 268714 800
rect 269210 0 269266 800
rect 269854 0 269910 800
rect 270406 0 270462 800
rect 271050 0 271106 800
rect 271694 0 271750 800
rect 272246 0 272302 800
rect 272890 0 272946 800
rect 273442 0 273498 800
rect 274086 0 274142 800
rect 274730 0 274786 800
rect 275282 0 275338 800
rect 275926 0 275982 800
rect 276570 0 276626 800
rect 277122 0 277178 800
rect 277766 0 277822 800
rect 278318 0 278374 800
rect 278962 0 279018 800
rect 279606 0 279662 800
rect 280158 0 280214 800
rect 280802 0 280858 800
rect 281354 0 281410 800
rect 281998 0 282054 800
rect 282642 0 282698 800
rect 283194 0 283250 800
rect 283838 0 283894 800
rect 284482 0 284538 800
rect 285034 0 285090 800
rect 285678 0 285734 800
rect 286230 0 286286 800
rect 286874 0 286930 800
rect 287518 0 287574 800
rect 288070 0 288126 800
rect 288714 0 288770 800
rect 289266 0 289322 800
rect 289910 0 289966 800
rect 290554 0 290610 800
rect 291106 0 291162 800
rect 291750 0 291806 800
rect 292394 0 292450 800
rect 292946 0 293002 800
rect 293590 0 293646 800
rect 294142 0 294198 800
rect 294786 0 294842 800
rect 295430 0 295486 800
rect 295982 0 296038 800
rect 296626 0 296682 800
rect 297178 0 297234 800
rect 297822 0 297878 800
rect 298466 0 298522 800
rect 299018 0 299074 800
rect 299662 0 299718 800
<< obsm2 >>
rect 296 179144 1250 179200
rect 1418 179144 3826 179200
rect 3994 179144 6494 179200
rect 6662 179144 9070 179200
rect 9238 179144 11738 179200
rect 11906 179144 14406 179200
rect 14574 179144 16982 179200
rect 17150 179144 19650 179200
rect 19818 179144 22226 179200
rect 22394 179144 24894 179200
rect 25062 179144 27562 179200
rect 27730 179144 30138 179200
rect 30306 179144 32806 179200
rect 32974 179144 35382 179200
rect 35550 179144 38050 179200
rect 38218 179144 40718 179200
rect 40886 179144 43294 179200
rect 43462 179144 45962 179200
rect 46130 179144 48538 179200
rect 48706 179144 51206 179200
rect 51374 179144 53874 179200
rect 54042 179144 56450 179200
rect 56618 179144 59118 179200
rect 59286 179144 61694 179200
rect 61862 179144 64362 179200
rect 64530 179144 67030 179200
rect 67198 179144 69606 179200
rect 69774 179144 72274 179200
rect 72442 179144 74850 179200
rect 75018 179144 77518 179200
rect 77686 179144 80186 179200
rect 80354 179144 82762 179200
rect 82930 179144 85430 179200
rect 85598 179144 88006 179200
rect 88174 179144 90674 179200
rect 90842 179144 93342 179200
rect 93510 179144 95918 179200
rect 96086 179144 98586 179200
rect 98754 179144 101254 179200
rect 101422 179144 103830 179200
rect 103998 179144 106498 179200
rect 106666 179144 109074 179200
rect 109242 179144 111742 179200
rect 111910 179144 114410 179200
rect 114578 179144 116986 179200
rect 117154 179144 119654 179200
rect 119822 179144 122230 179200
rect 122398 179144 124898 179200
rect 125066 179144 127566 179200
rect 127734 179144 130142 179200
rect 130310 179144 132810 179200
rect 132978 179144 135386 179200
rect 135554 179144 138054 179200
rect 138222 179144 140722 179200
rect 140890 179144 143298 179200
rect 143466 179144 145966 179200
rect 146134 179144 148542 179200
rect 148710 179144 151210 179200
rect 151378 179144 153878 179200
rect 154046 179144 156454 179200
rect 156622 179144 159122 179200
rect 159290 179144 161698 179200
rect 161866 179144 164366 179200
rect 164534 179144 167034 179200
rect 167202 179144 169610 179200
rect 169778 179144 172278 179200
rect 172446 179144 174854 179200
rect 175022 179144 177522 179200
rect 177690 179144 180190 179200
rect 180358 179144 182766 179200
rect 182934 179144 185434 179200
rect 185602 179144 188010 179200
rect 188178 179144 190678 179200
rect 190846 179144 193346 179200
rect 193514 179144 195922 179200
rect 196090 179144 198590 179200
rect 198758 179144 201258 179200
rect 201426 179144 203834 179200
rect 204002 179144 206502 179200
rect 206670 179144 209078 179200
rect 209246 179144 211746 179200
rect 211914 179144 214414 179200
rect 214582 179144 216990 179200
rect 217158 179144 219658 179200
rect 219826 179144 222234 179200
rect 222402 179144 224902 179200
rect 225070 179144 227570 179200
rect 227738 179144 230146 179200
rect 230314 179144 232814 179200
rect 232982 179144 235390 179200
rect 235558 179144 238058 179200
rect 238226 179144 240726 179200
rect 240894 179144 243302 179200
rect 243470 179144 245970 179200
rect 246138 179144 248546 179200
rect 248714 179144 251214 179200
rect 251382 179144 253882 179200
rect 254050 179144 256458 179200
rect 256626 179144 259126 179200
rect 259294 179144 261702 179200
rect 261870 179144 264370 179200
rect 264538 179144 267038 179200
rect 267206 179144 269614 179200
rect 269782 179144 272282 179200
rect 272450 179144 274858 179200
rect 275026 179144 277526 179200
rect 277694 179144 280194 179200
rect 280362 179144 282770 179200
rect 282938 179144 285438 179200
rect 285606 179144 288014 179200
rect 288182 179144 290682 179200
rect 290850 179144 293350 179200
rect 293518 179144 295926 179200
rect 296094 179144 298594 179200
rect 298762 179144 299716 179200
rect 296 856 299716 179144
rect 406 734 790 856
rect 958 734 1434 856
rect 1602 734 1986 856
rect 2154 734 2630 856
rect 2798 734 3274 856
rect 3442 734 3826 856
rect 3994 734 4470 856
rect 4638 734 5022 856
rect 5190 734 5666 856
rect 5834 734 6310 856
rect 6478 734 6862 856
rect 7030 734 7506 856
rect 7674 734 8058 856
rect 8226 734 8702 856
rect 8870 734 9346 856
rect 9514 734 9898 856
rect 10066 734 10542 856
rect 10710 734 11186 856
rect 11354 734 11738 856
rect 11906 734 12382 856
rect 12550 734 12934 856
rect 13102 734 13578 856
rect 13746 734 14222 856
rect 14390 734 14774 856
rect 14942 734 15418 856
rect 15586 734 15970 856
rect 16138 734 16614 856
rect 16782 734 17258 856
rect 17426 734 17810 856
rect 17978 734 18454 856
rect 18622 734 19098 856
rect 19266 734 19650 856
rect 19818 734 20294 856
rect 20462 734 20846 856
rect 21014 734 21490 856
rect 21658 734 22134 856
rect 22302 734 22686 856
rect 22854 734 23330 856
rect 23498 734 23882 856
rect 24050 734 24526 856
rect 24694 734 25170 856
rect 25338 734 25722 856
rect 25890 734 26366 856
rect 26534 734 27010 856
rect 27178 734 27562 856
rect 27730 734 28206 856
rect 28374 734 28758 856
rect 28926 734 29402 856
rect 29570 734 30046 856
rect 30214 734 30598 856
rect 30766 734 31242 856
rect 31410 734 31794 856
rect 31962 734 32438 856
rect 32606 734 33082 856
rect 33250 734 33634 856
rect 33802 734 34278 856
rect 34446 734 34922 856
rect 35090 734 35474 856
rect 35642 734 36118 856
rect 36286 734 36670 856
rect 36838 734 37314 856
rect 37482 734 37958 856
rect 38126 734 38510 856
rect 38678 734 39154 856
rect 39322 734 39706 856
rect 39874 734 40350 856
rect 40518 734 40994 856
rect 41162 734 41546 856
rect 41714 734 42190 856
rect 42358 734 42834 856
rect 43002 734 43386 856
rect 43554 734 44030 856
rect 44198 734 44582 856
rect 44750 734 45226 856
rect 45394 734 45870 856
rect 46038 734 46422 856
rect 46590 734 47066 856
rect 47234 734 47618 856
rect 47786 734 48262 856
rect 48430 734 48906 856
rect 49074 734 49458 856
rect 49626 734 50102 856
rect 50270 734 50746 856
rect 50914 734 51298 856
rect 51466 734 51942 856
rect 52110 734 52494 856
rect 52662 734 53138 856
rect 53306 734 53782 856
rect 53950 734 54334 856
rect 54502 734 54978 856
rect 55146 734 55530 856
rect 55698 734 56174 856
rect 56342 734 56818 856
rect 56986 734 57370 856
rect 57538 734 58014 856
rect 58182 734 58658 856
rect 58826 734 59210 856
rect 59378 734 59854 856
rect 60022 734 60406 856
rect 60574 734 61050 856
rect 61218 734 61694 856
rect 61862 734 62246 856
rect 62414 734 62890 856
rect 63058 734 63442 856
rect 63610 734 64086 856
rect 64254 734 64730 856
rect 64898 734 65282 856
rect 65450 734 65926 856
rect 66094 734 66478 856
rect 66646 734 67122 856
rect 67290 734 67766 856
rect 67934 734 68318 856
rect 68486 734 68962 856
rect 69130 734 69606 856
rect 69774 734 70158 856
rect 70326 734 70802 856
rect 70970 734 71354 856
rect 71522 734 71998 856
rect 72166 734 72642 856
rect 72810 734 73194 856
rect 73362 734 73838 856
rect 74006 734 74390 856
rect 74558 734 75034 856
rect 75202 734 75678 856
rect 75846 734 76230 856
rect 76398 734 76874 856
rect 77042 734 77518 856
rect 77686 734 78070 856
rect 78238 734 78714 856
rect 78882 734 79266 856
rect 79434 734 79910 856
rect 80078 734 80554 856
rect 80722 734 81106 856
rect 81274 734 81750 856
rect 81918 734 82302 856
rect 82470 734 82946 856
rect 83114 734 83590 856
rect 83758 734 84142 856
rect 84310 734 84786 856
rect 84954 734 85430 856
rect 85598 734 85982 856
rect 86150 734 86626 856
rect 86794 734 87178 856
rect 87346 734 87822 856
rect 87990 734 88466 856
rect 88634 734 89018 856
rect 89186 734 89662 856
rect 89830 734 90214 856
rect 90382 734 90858 856
rect 91026 734 91502 856
rect 91670 734 92054 856
rect 92222 734 92698 856
rect 92866 734 93342 856
rect 93510 734 93894 856
rect 94062 734 94538 856
rect 94706 734 95090 856
rect 95258 734 95734 856
rect 95902 734 96378 856
rect 96546 734 96930 856
rect 97098 734 97574 856
rect 97742 734 98126 856
rect 98294 734 98770 856
rect 98938 734 99414 856
rect 99582 734 99966 856
rect 100134 734 100610 856
rect 100778 734 101254 856
rect 101422 734 101806 856
rect 101974 734 102450 856
rect 102618 734 103002 856
rect 103170 734 103646 856
rect 103814 734 104290 856
rect 104458 734 104842 856
rect 105010 734 105486 856
rect 105654 734 106038 856
rect 106206 734 106682 856
rect 106850 734 107326 856
rect 107494 734 107878 856
rect 108046 734 108522 856
rect 108690 734 109166 856
rect 109334 734 109718 856
rect 109886 734 110362 856
rect 110530 734 110914 856
rect 111082 734 111558 856
rect 111726 734 112202 856
rect 112370 734 112754 856
rect 112922 734 113398 856
rect 113566 734 113950 856
rect 114118 734 114594 856
rect 114762 734 115238 856
rect 115406 734 115790 856
rect 115958 734 116434 856
rect 116602 734 117078 856
rect 117246 734 117630 856
rect 117798 734 118274 856
rect 118442 734 118826 856
rect 118994 734 119470 856
rect 119638 734 120114 856
rect 120282 734 120666 856
rect 120834 734 121310 856
rect 121478 734 121862 856
rect 122030 734 122506 856
rect 122674 734 123150 856
rect 123318 734 123702 856
rect 123870 734 124346 856
rect 124514 734 124898 856
rect 125066 734 125542 856
rect 125710 734 126186 856
rect 126354 734 126738 856
rect 126906 734 127382 856
rect 127550 734 128026 856
rect 128194 734 128578 856
rect 128746 734 129222 856
rect 129390 734 129774 856
rect 129942 734 130418 856
rect 130586 734 131062 856
rect 131230 734 131614 856
rect 131782 734 132258 856
rect 132426 734 132810 856
rect 132978 734 133454 856
rect 133622 734 134098 856
rect 134266 734 134650 856
rect 134818 734 135294 856
rect 135462 734 135938 856
rect 136106 734 136490 856
rect 136658 734 137134 856
rect 137302 734 137686 856
rect 137854 734 138330 856
rect 138498 734 138974 856
rect 139142 734 139526 856
rect 139694 734 140170 856
rect 140338 734 140722 856
rect 140890 734 141366 856
rect 141534 734 142010 856
rect 142178 734 142562 856
rect 142730 734 143206 856
rect 143374 734 143850 856
rect 144018 734 144402 856
rect 144570 734 145046 856
rect 145214 734 145598 856
rect 145766 734 146242 856
rect 146410 734 146886 856
rect 147054 734 147438 856
rect 147606 734 148082 856
rect 148250 734 148634 856
rect 148802 734 149278 856
rect 149446 734 149922 856
rect 150090 734 150474 856
rect 150642 734 151118 856
rect 151286 734 151762 856
rect 151930 734 152314 856
rect 152482 734 152958 856
rect 153126 734 153510 856
rect 153678 734 154154 856
rect 154322 734 154798 856
rect 154966 734 155350 856
rect 155518 734 155994 856
rect 156162 734 156546 856
rect 156714 734 157190 856
rect 157358 734 157834 856
rect 158002 734 158386 856
rect 158554 734 159030 856
rect 159198 734 159674 856
rect 159842 734 160226 856
rect 160394 734 160870 856
rect 161038 734 161422 856
rect 161590 734 162066 856
rect 162234 734 162710 856
rect 162878 734 163262 856
rect 163430 734 163906 856
rect 164074 734 164458 856
rect 164626 734 165102 856
rect 165270 734 165746 856
rect 165914 734 166298 856
rect 166466 734 166942 856
rect 167110 734 167586 856
rect 167754 734 168138 856
rect 168306 734 168782 856
rect 168950 734 169334 856
rect 169502 734 169978 856
rect 170146 734 170622 856
rect 170790 734 171174 856
rect 171342 734 171818 856
rect 171986 734 172370 856
rect 172538 734 173014 856
rect 173182 734 173658 856
rect 173826 734 174210 856
rect 174378 734 174854 856
rect 175022 734 175498 856
rect 175666 734 176050 856
rect 176218 734 176694 856
rect 176862 734 177246 856
rect 177414 734 177890 856
rect 178058 734 178534 856
rect 178702 734 179086 856
rect 179254 734 179730 856
rect 179898 734 180282 856
rect 180450 734 180926 856
rect 181094 734 181570 856
rect 181738 734 182122 856
rect 182290 734 182766 856
rect 182934 734 183318 856
rect 183486 734 183962 856
rect 184130 734 184606 856
rect 184774 734 185158 856
rect 185326 734 185802 856
rect 185970 734 186446 856
rect 186614 734 186998 856
rect 187166 734 187642 856
rect 187810 734 188194 856
rect 188362 734 188838 856
rect 189006 734 189482 856
rect 189650 734 190034 856
rect 190202 734 190678 856
rect 190846 734 191230 856
rect 191398 734 191874 856
rect 192042 734 192518 856
rect 192686 734 193070 856
rect 193238 734 193714 856
rect 193882 734 194358 856
rect 194526 734 194910 856
rect 195078 734 195554 856
rect 195722 734 196106 856
rect 196274 734 196750 856
rect 196918 734 197394 856
rect 197562 734 197946 856
rect 198114 734 198590 856
rect 198758 734 199142 856
rect 199310 734 199786 856
rect 199954 734 200430 856
rect 200598 734 200982 856
rect 201150 734 201626 856
rect 201794 734 202270 856
rect 202438 734 202822 856
rect 202990 734 203466 856
rect 203634 734 204018 856
rect 204186 734 204662 856
rect 204830 734 205306 856
rect 205474 734 205858 856
rect 206026 734 206502 856
rect 206670 734 207054 856
rect 207222 734 207698 856
rect 207866 734 208342 856
rect 208510 734 208894 856
rect 209062 734 209538 856
rect 209706 734 210182 856
rect 210350 734 210734 856
rect 210902 734 211378 856
rect 211546 734 211930 856
rect 212098 734 212574 856
rect 212742 734 213218 856
rect 213386 734 213770 856
rect 213938 734 214414 856
rect 214582 734 214966 856
rect 215134 734 215610 856
rect 215778 734 216254 856
rect 216422 734 216806 856
rect 216974 734 217450 856
rect 217618 734 218094 856
rect 218262 734 218646 856
rect 218814 734 219290 856
rect 219458 734 219842 856
rect 220010 734 220486 856
rect 220654 734 221130 856
rect 221298 734 221682 856
rect 221850 734 222326 856
rect 222494 734 222878 856
rect 223046 734 223522 856
rect 223690 734 224166 856
rect 224334 734 224718 856
rect 224886 734 225362 856
rect 225530 734 226006 856
rect 226174 734 226558 856
rect 226726 734 227202 856
rect 227370 734 227754 856
rect 227922 734 228398 856
rect 228566 734 229042 856
rect 229210 734 229594 856
rect 229762 734 230238 856
rect 230406 734 230790 856
rect 230958 734 231434 856
rect 231602 734 232078 856
rect 232246 734 232630 856
rect 232798 734 233274 856
rect 233442 734 233918 856
rect 234086 734 234470 856
rect 234638 734 235114 856
rect 235282 734 235666 856
rect 235834 734 236310 856
rect 236478 734 236954 856
rect 237122 734 237506 856
rect 237674 734 238150 856
rect 238318 734 238702 856
rect 238870 734 239346 856
rect 239514 734 239990 856
rect 240158 734 240542 856
rect 240710 734 241186 856
rect 241354 734 241738 856
rect 241906 734 242382 856
rect 242550 734 243026 856
rect 243194 734 243578 856
rect 243746 734 244222 856
rect 244390 734 244866 856
rect 245034 734 245418 856
rect 245586 734 246062 856
rect 246230 734 246614 856
rect 246782 734 247258 856
rect 247426 734 247902 856
rect 248070 734 248454 856
rect 248622 734 249098 856
rect 249266 734 249650 856
rect 249818 734 250294 856
rect 250462 734 250938 856
rect 251106 734 251490 856
rect 251658 734 252134 856
rect 252302 734 252778 856
rect 252946 734 253330 856
rect 253498 734 253974 856
rect 254142 734 254526 856
rect 254694 734 255170 856
rect 255338 734 255814 856
rect 255982 734 256366 856
rect 256534 734 257010 856
rect 257178 734 257562 856
rect 257730 734 258206 856
rect 258374 734 258850 856
rect 259018 734 259402 856
rect 259570 734 260046 856
rect 260214 734 260690 856
rect 260858 734 261242 856
rect 261410 734 261886 856
rect 262054 734 262438 856
rect 262606 734 263082 856
rect 263250 734 263726 856
rect 263894 734 264278 856
rect 264446 734 264922 856
rect 265090 734 265474 856
rect 265642 734 266118 856
rect 266286 734 266762 856
rect 266930 734 267314 856
rect 267482 734 267958 856
rect 268126 734 268602 856
rect 268770 734 269154 856
rect 269322 734 269798 856
rect 269966 734 270350 856
rect 270518 734 270994 856
rect 271162 734 271638 856
rect 271806 734 272190 856
rect 272358 734 272834 856
rect 273002 734 273386 856
rect 273554 734 274030 856
rect 274198 734 274674 856
rect 274842 734 275226 856
rect 275394 734 275870 856
rect 276038 734 276514 856
rect 276682 734 277066 856
rect 277234 734 277710 856
rect 277878 734 278262 856
rect 278430 734 278906 856
rect 279074 734 279550 856
rect 279718 734 280102 856
rect 280270 734 280746 856
rect 280914 734 281298 856
rect 281466 734 281942 856
rect 282110 734 282586 856
rect 282754 734 283138 856
rect 283306 734 283782 856
rect 283950 734 284426 856
rect 284594 734 284978 856
rect 285146 734 285622 856
rect 285790 734 286174 856
rect 286342 734 286818 856
rect 286986 734 287462 856
rect 287630 734 288014 856
rect 288182 734 288658 856
rect 288826 734 289210 856
rect 289378 734 289854 856
rect 290022 734 290498 856
rect 290666 734 291050 856
rect 291218 734 291694 856
rect 291862 734 292338 856
rect 292506 734 292890 856
rect 293058 734 293534 856
rect 293702 734 294086 856
rect 294254 734 294730 856
rect 294898 734 295374 856
rect 295542 734 295926 856
rect 296094 734 296570 856
rect 296738 734 297122 856
rect 297290 734 297766 856
rect 297934 734 298410 856
rect 298578 734 298962 856
rect 299130 734 299606 856
<< metal3 >>
rect 299200 90040 300000 90160
<< obsm3 >>
rect 1301 2143 296368 177377
<< metal4 >>
rect 4208 2128 4528 177392
rect 19568 2128 19888 177392
rect 34928 2128 35248 177392
rect 50288 2128 50608 177392
rect 65648 2128 65968 177392
rect 81008 2128 81328 177392
rect 96368 2128 96688 177392
rect 111728 2128 112048 177392
rect 127088 2128 127408 177392
rect 142448 2128 142768 177392
rect 157808 2128 158128 177392
rect 173168 2128 173488 177392
rect 188528 2128 188848 177392
rect 203888 2128 204208 177392
rect 219248 2128 219568 177392
rect 234608 2128 234928 177392
rect 249968 2128 250288 177392
rect 265328 2128 265648 177392
rect 280688 2128 281008 177392
rect 296048 2128 296368 177392
<< obsm4 >>
rect 34467 54843 34848 154597
rect 35328 54843 50208 154597
rect 50688 54843 65568 154597
rect 66048 54843 80928 154597
rect 81408 54843 96288 154597
rect 96768 54843 111648 154597
rect 112128 54843 127008 154597
rect 127488 54843 142368 154597
rect 142848 54843 149901 154597
<< labels >>
rlabel metal2 s 1306 179200 1362 180000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 80242 179200 80298 180000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 88062 179200 88118 180000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 95974 179200 96030 180000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 103886 179200 103942 180000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 111798 179200 111854 180000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 119710 179200 119766 180000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 127622 179200 127678 180000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 135442 179200 135498 180000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 143354 179200 143410 180000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 151266 179200 151322 180000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 9126 179200 9182 180000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 159178 179200 159234 180000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 167090 179200 167146 180000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 174910 179200 174966 180000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 182822 179200 182878 180000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 190734 179200 190790 180000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 198646 179200 198702 180000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 206558 179200 206614 180000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 214470 179200 214526 180000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 222290 179200 222346 180000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 230202 179200 230258 180000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 17038 179200 17094 180000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 238114 179200 238170 180000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 246026 179200 246082 180000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 253938 179200 253994 180000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 261758 179200 261814 180000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 269670 179200 269726 180000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 277582 179200 277638 180000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 285494 179200 285550 180000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 293406 179200 293462 180000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 24950 179200 25006 180000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 32862 179200 32918 180000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 40774 179200 40830 180000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 48594 179200 48650 180000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 56506 179200 56562 180000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 64418 179200 64474 180000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 72330 179200 72386 180000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3882 179200 3938 180000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 82818 179200 82874 180000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 90730 179200 90786 180000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 98642 179200 98698 180000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 106554 179200 106610 180000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 114466 179200 114522 180000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 122286 179200 122342 180000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 130198 179200 130254 180000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 138110 179200 138166 180000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 146022 179200 146078 180000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 153934 179200 153990 180000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 11794 179200 11850 180000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 161754 179200 161810 180000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 169666 179200 169722 180000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 177578 179200 177634 180000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 185490 179200 185546 180000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 193402 179200 193458 180000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 201314 179200 201370 180000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 209134 179200 209190 180000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 217046 179200 217102 180000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 224958 179200 225014 180000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 232870 179200 232926 180000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 19706 179200 19762 180000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 240782 179200 240838 180000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 248602 179200 248658 180000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 256514 179200 256570 180000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 264426 179200 264482 180000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 272338 179200 272394 180000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 280250 179200 280306 180000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 288070 179200 288126 180000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 295982 179200 296038 180000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 27618 179200 27674 180000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 35438 179200 35494 180000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 43350 179200 43406 180000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 51262 179200 51318 180000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 59174 179200 59230 180000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 67086 179200 67142 180000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 74906 179200 74962 180000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 6550 179200 6606 180000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 85486 179200 85542 180000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 93398 179200 93454 180000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 101310 179200 101366 180000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 109130 179200 109186 180000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 117042 179200 117098 180000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 124954 179200 125010 180000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 132866 179200 132922 180000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 140778 179200 140834 180000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 148598 179200 148654 180000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 156510 179200 156566 180000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 14462 179200 14518 180000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 164422 179200 164478 180000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 172334 179200 172390 180000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 180246 179200 180302 180000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 188066 179200 188122 180000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 195978 179200 196034 180000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 203890 179200 203946 180000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 211802 179200 211858 180000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 219714 179200 219770 180000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 227626 179200 227682 180000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 235446 179200 235502 180000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 22282 179200 22338 180000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 243358 179200 243414 180000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 251270 179200 251326 180000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 259182 179200 259238 180000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 267094 179200 267150 180000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 274914 179200 274970 180000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 282826 179200 282882 180000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 290738 179200 290794 180000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 298650 179200 298706 180000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 30194 179200 30250 180000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 38106 179200 38162 180000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 46018 179200 46074 180000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 53930 179200 53986 180000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 61750 179200 61806 180000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 69662 179200 69718 180000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 77574 179200 77630 180000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 298466 0 298522 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 299018 0 299074 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 299662 0 299718 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 247314 0 247370 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 249154 0 249210 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 250994 0 251050 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 252834 0 252890 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 254582 0 254638 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 256422 0 256478 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 258262 0 258318 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 260102 0 260158 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 261942 0 261998 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 263782 0 263838 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 265530 0 265586 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 267370 0 267426 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 269210 0 269266 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 271050 0 271106 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 272890 0 272946 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 274730 0 274786 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 276570 0 276626 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 278318 0 278374 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 280158 0 280214 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 281998 0 282054 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 283838 0 283894 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 285678 0 285734 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 287518 0 287574 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 289266 0 289322 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 291106 0 291162 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 292946 0 293002 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 294786 0 294842 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 296626 0 296682 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 123206 0 123262 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 128634 0 128690 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 134154 0 134210 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 137742 0 137798 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 139582 0 139638 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 141422 0 141478 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 143262 0 143318 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 150530 0 150586 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 152370 0 152426 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 154210 0 154266 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 156050 0 156106 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 157890 0 157946 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 161478 0 161534 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 163318 0 163374 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 165158 0 165214 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 166998 0 167054 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 168838 0 168894 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 170678 0 170734 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 172426 0 172482 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 177946 0 178002 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 179786 0 179842 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 181626 0 181682 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 183374 0 183430 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 185214 0 185270 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 187054 0 187110 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 188894 0 188950 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 190734 0 190790 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 192574 0 192630 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 194414 0 194470 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 196162 0 196218 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 198002 0 198058 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 199842 0 199898 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 201682 0 201738 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 203522 0 203578 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 205362 0 205418 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 207110 0 207166 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 208950 0 209006 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 210790 0 210846 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 212630 0 212686 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 214470 0 214526 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 216310 0 216366 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 218150 0 218206 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 219898 0 219954 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 221738 0 221794 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 223578 0 223634 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 225418 0 225474 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 227258 0 227314 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 229098 0 229154 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 230846 0 230902 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 232686 0 232742 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 234526 0 234582 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 236366 0 236422 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 238206 0 238262 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 240046 0 240102 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 241794 0 241850 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 243634 0 243690 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 245474 0 245530 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 247958 0 248014 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 249706 0 249762 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 251546 0 251602 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 253386 0 253442 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 255226 0 255282 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 257066 0 257122 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 258906 0 258962 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 260746 0 260802 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 262494 0 262550 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 264334 0 264390 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 266174 0 266230 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 268014 0 268070 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 269854 0 269910 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 271694 0 271750 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 273442 0 273498 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 275282 0 275338 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 277122 0 277178 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 278962 0 279018 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 280802 0 280858 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 282642 0 282698 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 85486 0 85542 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 284482 0 284538 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 286230 0 286286 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 288070 0 288126 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 289910 0 289966 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 291750 0 291806 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 293590 0 293646 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 295430 0 295486 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 297178 0 297234 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 89074 0 89130 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 90914 0 90970 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 94594 0 94650 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 96434 0 96490 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 98182 0 98238 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 100022 0 100078 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 101862 0 101918 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 103702 0 103758 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 107382 0 107438 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 110970 0 111026 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 112810 0 112866 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 116490 0 116546 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 118330 0 118386 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 120170 0 120226 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 127438 0 127494 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 129278 0 129334 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 131118 0 131174 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 132866 0 132922 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 134706 0 134762 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 136546 0 136602 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 138386 0 138442 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 140226 0 140282 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 142066 0 142122 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 143906 0 143962 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 145654 0 145710 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 147494 0 147550 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 149334 0 149390 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 151174 0 151230 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 153014 0 153070 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 154854 0 154910 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 156602 0 156658 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 158442 0 158498 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 160282 0 160338 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 162122 0 162178 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 163962 0 164018 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 165802 0 165858 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 167642 0 167698 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 169390 0 169446 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 171230 0 171286 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 173070 0 173126 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 174910 0 174966 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 176750 0 176806 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 178590 0 178646 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 180338 0 180394 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 182178 0 182234 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 184018 0 184074 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 185858 0 185914 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 187698 0 187754 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 189538 0 189594 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 191286 0 191342 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 76286 0 76342 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 193126 0 193182 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 194966 0 195022 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 196806 0 196862 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 198646 0 198702 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 200486 0 200542 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 202326 0 202382 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 204074 0 204130 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 205914 0 205970 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 207754 0 207810 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 209594 0 209650 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 211434 0 211490 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 213274 0 213330 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 215022 0 215078 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 216862 0 216918 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 218702 0 218758 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 220542 0 220598 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 222382 0 222438 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 224222 0 224278 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 226062 0 226118 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 227810 0 227866 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 79966 0 80022 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 229650 0 229706 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 231490 0 231546 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 233330 0 233386 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 235170 0 235226 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 237010 0 237066 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 238758 0 238814 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 240598 0 240654 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 242438 0 242494 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 244278 0 244334 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 246118 0 246174 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 65982 0 66038 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 248510 0 248566 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 250350 0 250406 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 252190 0 252246 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 254030 0 254086 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 255870 0 255926 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 257618 0 257674 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 259458 0 259514 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 261298 0 261354 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 263138 0 263194 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 264978 0 265034 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 266818 0 266874 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 268658 0 268714 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 270406 0 270462 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 272246 0 272302 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 274086 0 274142 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 275926 0 275982 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 277766 0 277822 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 279606 0 279662 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 281354 0 281410 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 283194 0 283250 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 285034 0 285090 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 286874 0 286930 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 288714 0 288770 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 290554 0 290610 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 292394 0 292450 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 294142 0 294198 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 295982 0 296038 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 297822 0 297878 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 129830 0 129886 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 131670 0 131726 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 137190 0 137246 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 139030 0 139086 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 140778 0 140834 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 151818 0 151874 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 157246 0 157302 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 159086 0 159142 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 160926 0 160982 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 164514 0 164570 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 166354 0 166410 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 168194 0 168250 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 170034 0 170090 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 171874 0 171930 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 173714 0 173770 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 175554 0 175610 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 177302 0 177358 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 179142 0 179198 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 182822 0 182878 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 184662 0 184718 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 186502 0 186558 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 188250 0 188306 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 190090 0 190146 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 191930 0 191986 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 193770 0 193826 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 195610 0 195666 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 197450 0 197506 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 199198 0 199254 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 201038 0 201094 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 202878 0 202934 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 204718 0 204774 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 206558 0 206614 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 208398 0 208454 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 210238 0 210294 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 211986 0 212042 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 213826 0 213882 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 215666 0 215722 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 217506 0 217562 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 219346 0 219402 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 221186 0 221242 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 222934 0 222990 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 224774 0 224830 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 226614 0 226670 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 228454 0 228510 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 230294 0 230350 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 232134 0 232190 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 233974 0 234030 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 235722 0 235778 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 237562 0 237618 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 239402 0 239458 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 241242 0 241298 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 243082 0 243138 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 244922 0 244978 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 246670 0 246726 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal3 s 299200 90040 300000 90160 6 user_clock2
port 502 nsew signal input
rlabel metal4 s 4208 2128 4528 177392 6 vccd1
port 503 nsew power input
rlabel metal4 s 34928 2128 35248 177392 6 vccd1
port 503 nsew power input
rlabel metal4 s 65648 2128 65968 177392 6 vccd1
port 503 nsew power input
rlabel metal4 s 96368 2128 96688 177392 6 vccd1
port 503 nsew power input
rlabel metal4 s 127088 2128 127408 177392 6 vccd1
port 503 nsew power input
rlabel metal4 s 157808 2128 158128 177392 6 vccd1
port 503 nsew power input
rlabel metal4 s 188528 2128 188848 177392 6 vccd1
port 503 nsew power input
rlabel metal4 s 219248 2128 219568 177392 6 vccd1
port 503 nsew power input
rlabel metal4 s 249968 2128 250288 177392 6 vccd1
port 503 nsew power input
rlabel metal4 s 280688 2128 281008 177392 6 vccd1
port 503 nsew power input
rlabel metal4 s 19568 2128 19888 177392 6 vssd1
port 504 nsew ground input
rlabel metal4 s 50288 2128 50608 177392 6 vssd1
port 504 nsew ground input
rlabel metal4 s 81008 2128 81328 177392 6 vssd1
port 504 nsew ground input
rlabel metal4 s 111728 2128 112048 177392 6 vssd1
port 504 nsew ground input
rlabel metal4 s 142448 2128 142768 177392 6 vssd1
port 504 nsew ground input
rlabel metal4 s 173168 2128 173488 177392 6 vssd1
port 504 nsew ground input
rlabel metal4 s 203888 2128 204208 177392 6 vssd1
port 504 nsew ground input
rlabel metal4 s 234608 2128 234928 177392 6 vssd1
port 504 nsew ground input
rlabel metal4 s 265328 2128 265648 177392 6 vssd1
port 504 nsew ground input
rlabel metal4 s 296048 2128 296368 177392 6 vssd1
port 504 nsew ground input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 505 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 506 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_ack_o
port 507 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 wbs_adr_i[0]
port 508 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[10]
port 509 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_adr_i[11]
port 510 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wbs_adr_i[12]
port 511 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_adr_i[13]
port 512 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_adr_i[14]
port 513 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_adr_i[15]
port 514 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wbs_adr_i[16]
port 515 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 wbs_adr_i[17]
port 516 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 wbs_adr_i[18]
port 517 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 wbs_adr_i[19]
port 518 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_adr_i[1]
port 519 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 wbs_adr_i[20]
port 520 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 wbs_adr_i[21]
port 521 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wbs_adr_i[22]
port 522 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_adr_i[23]
port 523 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 wbs_adr_i[24]
port 524 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 wbs_adr_i[25]
port 525 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 wbs_adr_i[26]
port 526 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 wbs_adr_i[27]
port 527 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 wbs_adr_i[28]
port 528 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 wbs_adr_i[29]
port 529 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[2]
port 530 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 wbs_adr_i[30]
port 531 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 wbs_adr_i[31]
port 532 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[3]
port 533 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_adr_i[4]
port 534 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_adr_i[5]
port 535 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_adr_i[6]
port 536 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[7]
port 537 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[8]
port 538 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_adr_i[9]
port 539 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_cyc_i
port 540 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_dat_i[0]
port 541 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_i[10]
port 542 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wbs_dat_i[11]
port 543 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_i[12]
port 544 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 wbs_dat_i[13]
port 545 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_dat_i[14]
port 546 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_i[15]
port 547 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 wbs_dat_i[16]
port 548 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_i[17]
port 549 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 wbs_dat_i[18]
port 550 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_i[19]
port 551 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_i[1]
port 552 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 wbs_dat_i[20]
port 553 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 wbs_dat_i[21]
port 554 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 wbs_dat_i[22]
port 555 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 wbs_dat_i[23]
port 556 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 wbs_dat_i[24]
port 557 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 wbs_dat_i[25]
port 558 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wbs_dat_i[26]
port 559 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 wbs_dat_i[27]
port 560 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 wbs_dat_i[28]
port 561 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 wbs_dat_i[29]
port 562 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_i[2]
port 563 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 wbs_dat_i[30]
port 564 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 wbs_dat_i[31]
port 565 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_i[3]
port 566 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_i[4]
port 567 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_dat_i[5]
port 568 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_dat_i[6]
port 569 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_i[7]
port 570 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_i[8]
port 571 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_i[9]
port 572 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_o[0]
port 573 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_o[10]
port 574 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_o[11]
port 575 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_o[12]
port 576 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 wbs_dat_o[13]
port 577 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 wbs_dat_o[14]
port 578 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 wbs_dat_o[15]
port 579 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 wbs_dat_o[16]
port 580 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 wbs_dat_o[17]
port 581 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 wbs_dat_o[18]
port 582 nsew signal output
rlabel metal2 s 42246 0 42302 800 6 wbs_dat_o[19]
port 583 nsew signal output
rlabel metal2 s 7562 0 7618 800 6 wbs_dat_o[1]
port 584 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 wbs_dat_o[20]
port 585 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 wbs_dat_o[21]
port 586 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 wbs_dat_o[22]
port 587 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 wbs_dat_o[23]
port 588 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 wbs_dat_o[24]
port 589 nsew signal output
rlabel metal2 s 53194 0 53250 800 6 wbs_dat_o[25]
port 590 nsew signal output
rlabel metal2 s 55034 0 55090 800 6 wbs_dat_o[26]
port 591 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 wbs_dat_o[27]
port 592 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 wbs_dat_o[28]
port 593 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 wbs_dat_o[29]
port 594 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[2]
port 595 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 wbs_dat_o[30]
port 596 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 wbs_dat_o[31]
port 597 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_o[3]
port 598 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[4]
port 599 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_o[5]
port 600 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_o[6]
port 601 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_o[7]
port 602 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_o[8]
port 603 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_o[9]
port 604 nsew signal output
rlabel metal2 s 5722 0 5778 800 6 wbs_sel_i[0]
port 605 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_sel_i[1]
port 606 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_sel_i[2]
port 607 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_sel_i[3]
port 608 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_stb_i
port 609 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_we_i
port 610 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 300000 180000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 79418514
string GDS_START 1317242
<< end >>

